module helloWorld();
  
  initial begin
  	$display("Hello World");
  end
    
endmodule